�� t �Thu May 02 13:56:45 2024
PvP
1
CheckMate
White win
 1.  6664___       5153___
 2.  4644___       5344P__
 3.  5724___       4445___
 4.  3755___       0103___
 5.  2451__#       