�� t�Tue Apr 30 12:19:35 2024
PvP
1
CheckMate
White win
 1.  4644___       3133___
 2.  4433P__       4142___
 3.  3342P__       5142P__
 4.  5713__+       3031___
 5.  1331Q_+       4031B__
 6.  3764___       1022___
 7.  1725___       2234___
 8.  2513___       3413N__
 9.  2624___       0102___
10.  2413N__       0213P__
11.  1614___       1112___
12.  0717___       0002___
13.  1715___       0200___
14.  1545___       0001___
15.  6442P_+       3130___
16.  4535__+       2031___
17.  4231B_#       