�� t �Wed May 01 01:29:59 2024
PvP
1
CheckMate
White win
 1.  4644___       5153___
 2.  5724___       5344P__
 3.  3755___       4445___
 4.  2451__#       