�� tMWed May 01 14:10:11 2024
PvP
1
Timeout
Black win
 1.  5654___       6052___
 2.  4756___       5264__+
 3.  5655___       3133___
 4.  0605___       3032___
 5.  2624___       3324P__
 6.  1614___       3233__+
 7.  5565___       6476P__
 8.  1413___       7657B_+
 9.  6556___       2075___
10.  0706___       7060___
11.  0607___       6163___
12.  5463P__       6063P__
13.  6664___       6364P__
14.  1725___       3336P__
15.  3747___       3647Q_+
16.  5655___       4725N_+
17.  5556___       1022___
18.  1312___       0112P__
19.  0504___       0004P__
20.  0705___       0405R__
