�� t�Tue Apr 30 13:10:12 2024
PvP
1
CheckMate
White win
 1.  5654___       4143___
 2.  5443P__       6052___
 3.  6755___       6163___
 4.  6664___       5072___
 5.  5775___       O-O____
 6.  O-O____       5264P__
 7.  4644___       5153___
 8.  3746___       5344P__
 9.  4644P__       7261___
10.  4464N__       5055N__
11.  5755R__       6143P__
12.  6463P_+       6070___
13.  5565___       3041___
14.  6360__#       