�� t�Tue Apr 30 23:11:47 2024
PvP
1
Timeout
Black win
 1.  2624___       3133___
 2.  2433P__       3033P__
 3.  3715___       3315Q__
 4.  0615Q__       2123___
 5.  1725___       2324___
 6.  1524P__       2042___
 7.  3635___       4224P__
 8.  3524B__       1022___
 9.  2533___       2214___
10.  3325___       1426__+
11.  4737___       2607R__
12.  2504___       0715___
13.  0425___       1523___
14.  4644___       2344P__
15.  2544N__       5153___
16.  4465___       6052___
17.  6553P__       5244___
18.  5365___       4456P_+
19.  3747___       6163___
20.  6544___       6364___
21.  4456N__       6465___
22.  7665P__       5072___
23.  5644___       7227B__
24.  4737___       2716P__
25.  3747___       7173___
