�� t �Thu May 02 23:09:23 2024
PvP
1
CheckMate
White win
 1.  4644___       5153___
 2.  5724___       5344P__
 3.  3755___       4445___
 4.  2451__#       